-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Mon Nov 17 19:04:55 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY sentido_sm IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        hor : IN STD_LOGIC := '0';
        ahor : IN STD_LOGIC := '0';
        sentido0 : OUT STD_LOGIC;
        sentido1 : OUT STD_LOGIC
    );
END sentido_sm;

ARCHITECTURE BEHAVIOR OF sentido_sm IS
    TYPE type_fstate IS (cima,baixo,esq,dir);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,hor,ahor)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= cima;
            sentido0 <= '0';
            sentido1 <= '0';
        ELSE
            sentido0 <= '0';
            sentido1 <= '0';
            CASE fstate IS
                WHEN cima =>
                    IF (((ahor = '1') AND NOT((hor = '1')))) THEN
                        reg_fstate <= esq;
                    ELSIF (((hor = '1') AND NOT((ahor = '1')))) THEN
                        reg_fstate <= dir;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= cima;
                    END IF;

                    sentido0 <= '0';

                    sentido1 <= '0';
                WHEN baixo =>
                    IF (((ahor = '1') AND NOT((hor = '1')))) THEN
                        reg_fstate <= dir;
                    ELSIF (((hor = '1') AND NOT((ahor = '1')))) THEN
                        reg_fstate <= esq;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= baixo;
                    END IF;

                    sentido0 <= '0';

                    sentido1 <= '1';
                WHEN esq =>
                    IF (((ahor = '1') AND NOT((hor = '1')))) THEN
                        reg_fstate <= baixo;
                    ELSIF (((hor = '1') AND NOT((ahor = '1')))) THEN
                        reg_fstate <= cima;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= esq;
                    END IF;

                    sentido0 <= '1';

                    sentido1 <= '1';
                WHEN dir =>
                    IF (((ahor = '1') AND NOT((hor = '1')))) THEN
                        reg_fstate <= cima;
                    ELSIF (((hor = '1') AND NOT((ahor = '1')))) THEN
                        reg_fstate <= baixo;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= dir;
                    END IF;

                    sentido0 <= '1';

                    sentido1 <= '0';
                WHEN OTHERS => 
                    sentido0 <= 'X';
                    sentido1 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
