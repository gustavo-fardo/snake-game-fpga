clk1hz_inst : clk1hz PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
