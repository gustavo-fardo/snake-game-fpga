sentido_inst : sentido PORT MAP (
		clock	 => clock_sig,
		updown	 => updown_sig,
		q	 => q_sig
	);
